module Trojan(
   input  wire [3:0] a, b, c, d, e,
   input  wire [1:0] mode,
   output wire [7:0] y
);
   wire [7:0] m1, m2, m3, m4;

   assign m1 = (a + b) * (c + d);
   assign m2 = (a * c) + (b * d);
   assign m3 = ((a ^ b) + d) * (e ^ 4'b1010);
   assign m4 = (m1 + m2) ^ (m3 >> 1);
   assign y = (mode == 2'b00) ? m1 :
              (mode == 2'b01) ? m4 :
              (mode == 2'b10) ? m2 : m3;

endmodule